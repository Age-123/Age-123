module blk (
  0_0_2,
  0_0_2_BL,
  64_0_2,
  64_0_2_BL,
  128_0_2,
  128_0_2_BL,
  0_0_3,
  0_0_3_BL,
  64_0_3,
  64_0_3_BL,
  128_0_3,
  128_0_3_BL,
  300_300_2,
  300_300_2_BL,
  364_300_2,
  364_300_2_BL,
  428_300_2,
  428_300_2_BL,
);
input 0_0_2_BL ;
input 64_0_2_BL ;
input 128_0_2_BL ;
input 0_0_3_BL ;
input 64_0_3_BL ;
input 128_0_3_BL ;
input 300_300_2_BL ;
input 364_300_2_BL ;
input 428_300_2_BL ;
output 0_0_2 ;
output 64_0_2 ;
output 128_0_2 ;
output 0_0_3 ;
output 64_0_3 ;
output 128_0_3 ;
output 300_300_2 ;
output 364_300_2 ;
output 428_300_2 ;
wire 0_0_2 ;
wire 0_0_2_BL ;
wire 64_0_2 ;
wire 64_0_2_BL ;
wire 128_0_2 ;
wire 128_0_2_BL ;
wire 0_0_3 ;
wire 0_0_3_BL ;
wire 64_0_3 ;
wire 64_0_3_BL ;
wire 128_0_3 ;
wire 128_0_3_BL ;
wire 300_300_2 ;
wire 300_300_2_BL ;
wire 364_300_2 ;
wire 364_300_2_BL ;
wire 428_300_2 ;
wire 428_300_2_BL ;
assign 0_0_2 = 0_0_2_BL ;
assign 64_0_2 = 64_0_2_BL ;
assign 128_0_2 = 128_0_2_BL ;
assign 0_0_3 = 0_0_3_BL ;
assign 64_0_3 = 64_0_3_BL ;
assign 128_0_3 = 128_0_3_BL ;
assign 300_300_2 = 300_300_2_BL ;
assign 364_300_2 = 364_300_2_BL ;
assign 428_300_2 = 428_300_2_BL ;
end module
